
`ifndef __UCSBIEEE__GPU__RTL__HEADERS__PARAMETERS_VH
`define __UCSBIEEE__GPU__RTL__HEADERS__PARAMETERS_VH


`define VRAM_SIZE       12'h900
`define VRAM_ADDR_WIDTH 12


`endif
