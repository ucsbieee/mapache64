
`define TEST_PMF    "vram-tests/random/pmf.dat"
`define TEST_PMB    "vram-tests/random/pmb.dat"
`define TEST_NTBL   "vram-tests/random/ntbl.dat"
`define TEST_OBM    "vram-tests/random/obm.dat"
