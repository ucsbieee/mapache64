
`ifndef __UCSBIEEE__TOP__SIM__HEADERS__TIMING_VH
`define __UCSBIEEE__TOP__SIM__HEADERS__TIMING_VH


`define TIMESCALE   1s/1fs

`define GPU_CLK_FREQ    12587500
`define GPU_CLK_PERIOD  ( 1.0 / `GPU_CLK_FREQ )

`endif
