
`define TIMESCALE   1s/1fs
