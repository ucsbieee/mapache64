
module clk_100_TO_clk_12_5875_m (
    output clk_12_5875,
    input clk_100
);

endmodule
