
struct {
    logic     [7:0] x       ;
    logic    [15:0] data    ;
    logic     [2:0] color   ;
    logic           valid   ;
} obsm[7:0];
