
`ifndef __UCSBIEEE__CONTROLLER_INTERFACE__SIM__TIMING_VH
`define __UCSBIEEE__CONTROLLER_INTERFACE__SIM__TIMING_VH


`define TIMESCALE   1s/1fs

`define CPU_CLK_FREQ    1000000
`define CPU_CLK_PERIOD  ( 1.0 / `CPU_CLK_FREQ )

`endif
