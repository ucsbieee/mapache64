
`define VRAM_SIZE       12'h900
`define VRAM_ADDR_WIDTH 12
