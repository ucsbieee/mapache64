
`define VRAM_SIZE       12'h900
`define VRAM_ADDR_WIDTH 12

`define GPU_CLK_FREQ    12587500
`define GPU_CLK_PERIOD  ( 1.0 / `GPU_CLK_FREQ )
